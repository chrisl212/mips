package mem_ftch_pkg;
  import mips_pkg::*;

  typedef struct packed {
    word_t      addr;
  } mem_ftch_pkt_t;
endpackage : mem_ftch_pkg
