package reg_file_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import reg_file_env_pkg::*;
  import reg_file_stim_pkg::*;

  `include "reg_file_test.svh"
endpackage : reg_file_tb_pkg
