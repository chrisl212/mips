package ftch_dec_pkg;
  typedef struct packed {
    word_t pc;
    word_t instr;
  } ftch_dec_pkt_t;
endpackage : ftch_dec_pkg
