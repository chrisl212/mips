typedef logic[`WORD_BITS-1:0] word_t;
