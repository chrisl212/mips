package cpu_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import cpu_env_pkg::*;
  import cpu_stim_pkg::*;

  `include "cpu_test.svh"
endpackage : cpu_tb_pkg
