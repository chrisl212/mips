package mem_env_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mips_pkg::*;
  import exec_mem_pkg::*;
  import mem_ftch_pkg::*;
  import mem_dmem_pkg::*;
  import mem_wrb_pkg::*;
  import haz_pkg::*;
  import clk_reset_iuvc_pkg::*;
  import exec_mem_iuvc_pkg::*;
  import mem_haz_iuvc_pkg::*;
  import mem_ftch_iuvc_pkg::*;
  import mem_dmem_iuvc_pkg::*;
  import dmem_mem_iuvc_pkg::*;
  import mem_wrb_iuvc_pkg::*;

  `include "mem_scoreboard.svh"
  `include "mem_env.svh"
endpackage : mem_env_pkg
