package reg_file_wr_req_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import reg_file_pkg::*;

  `include "reg_file_wr_req_seq_item.svh"
  `include "reg_file_wr_req_monitor.svh"
  `include "reg_file_wr_req_sequencer.svh"
  `include "reg_file_wr_req_master_driver.svh"
  `include "reg_file_wr_req_agent.svh"
endpackage : reg_file_wr_req_iuvc_pkg
