package instr_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mips_pkg::*;

  `include "instr.svh"
endpackage : instr_pkg
