package mem_ftch_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mem_ftch_pkg::*;

  `include "mem_ftch_seq_item.svh"
  `include "mem_ftch_monitor.svh"
  `include "mem_ftch_sequencer.svh"
  `include "mem_ftch_master_driver.svh"
  `include "mem_ftch_agent.svh"
endpackage : mem_ftch_iuvc_pkg
