package mem_stim_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mips_pkg::*;
  import clk_reset_iuvc_pkg::*;
  import exec_mem_iuvc_pkg::*;
  import mem_dmem_iuvc_pkg::*;
  import dmem_mem_iuvc_pkg::*;
  import mem_wrb_iuvc_pkg::*;

  `include "mem_virtual_sequencer.svh"
  `include "exec_mem_sequence.svh"
  `include "dmem_mem_sequence.svh"
  `include "mem_virtual_sequence.svh"
endpackage : mem_stim_pkg
