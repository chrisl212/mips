package alu_stim_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import alu_in_iuvc_pkg::*;
  import clk_reset_iuvc_pkg::*;

  `include "alu_virtual_sequencer.svh"
  `include "alu_in_sequence.svh"
  `include "alu_virtual_sequence.svh"
endpackage : alu_stim_pkg
