package ftch_imem_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import ftch_imem_pkg::*;

  `include "ftch_imem_seq_item.svh"
  `include "ftch_imem_monitor.svh"
  `include "ftch_imem_sequencer.svh"
  `include "ftch_imem_master_driver.svh"
  `include "ftch_imem_agent.svh"
endpackage : ftch_imem_iuvc_pkg
