package dec_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import dec_env_pkg::*;
  import dec_stim_pkg::*;

  `include "dec_test.svh"
endpackage : dec_tb_pkg
