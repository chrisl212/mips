package clk_reset_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "clk_reset_monitor.svh"
  `include "clk_reset_agent.svh"
endpackage : clk_reset_iuvc_pkg
