package alu_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import alu_env_pkg::*;
  import alu_stim_pkg::*;

  `include "alu_test.svh"
endpackage : alu_tb_pkg
