`define WORD_BITS (32)
