package exec_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import exec_env_pkg::*;
  import exec_stim_pkg::*;

  `include "exec_test.svh"
endpackage : exec_tb_pkg
