package imem_ftch_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import ftch_imem_pkg::*;

  `include "imem_ftch_seq_item.svh"
  `include "imem_ftch_monitor.svh"
  `include "imem_ftch_sequencer.svh"
  `include "imem_ftch_master_driver.svh"
  `include "imem_ftch_agent.svh"
endpackage : imem_ftch_iuvc_pkg
