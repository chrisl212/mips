package ftch_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import ftch_env_pkg::*;
  import ftch_stim_pkg::*;

  `include "ftch_test.svh"
endpackage : ftch_tb_pkg
