package mips_pkg;
  `include "common/defines.svh"
  `include "common/types.svh"
endpackage : mips_pkg

`include "intf/ftch_imem_pkg.svh"
`include "intf/ftch_dec_pkg.svh"
// `include "intf/dec_exec_pkg.svh"
// `include "intf/exec_mem_pkg.svh"
// `include "intf/mem_wrb_pkg.svh"
// `include "intf/wrb_dec_pkg.svh"
`include "intf/mem_ftch_pkg.svh"
`include "intf/reg_file_pkg.svh"
