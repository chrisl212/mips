package mem_tb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mem_env_pkg::*;
  import mem_stim_pkg::*;

  `include "mem_test.svh"
endpackage : mem_tb_pkg
