package ftch_env_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mips_pkg::*;
  import ftch_dec_pkg::*;
  import clk_reset_iuvc_pkg::*;
  import ftch_dec_iuvc_pkg::*;
  import ftch_imem_iuvc_pkg::*;
  import imem_ftch_iuvc_pkg::*;
  import mem_ftch_iuvc_pkg::*;

  `include "ftch_scoreboard.svh"
  `include "ftch_env.svh"
endpackage : ftch_env_pkg
