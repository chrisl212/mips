package mem_wrb_iuvc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import mem_wrb_pkg::*;
  
  `uvm_analysis_imp_decl(_mem_wrb)

  `include "mem_wrb_seq_item.svh"
  `include "mem_wrb_monitor.svh"
  `include "mem_wrb_sequencer.svh"
  `include "mem_wrb_master_driver.svh"
  `include "mem_wrb_agent.svh"
endpackage : mem_wrb_iuvc_pkg
